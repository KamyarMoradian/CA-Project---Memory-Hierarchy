library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
library work;
    use work.Types.ALL;

entity Processor is
    Port ( clk : in  STD_LOGIC;
           tlb_v : in  STD_LOGIC;
           cache_v : in  STD_LOGIC;
			  state_out : out state_type;
           data_out : out  STD_LOGIC_VECTOR (31 downto 0));
end Processor;

architecture Behavioral of Processor is

	-- =========================================================================
	-- Components:
	
	component Cache is
		Port ( read_en : in  STD_LOGIC;
				 write_en : in  STD_LOGIC;
             block_address : in  STD_LOGIC_VECTOR (10 downto 0); -- generated in Processor
             data_bus_in : in  STD_LOGIC_VECTOR (31 downto 0); -- coming from RAM
             clk : in  STD_LOGIC;
             hit : out  STD_LOGIC;
             data_bus_out : out  STD_LOGIC_VECTOR (31 downto 0));
	end component;

	component MainMemory is
		 Port ( read_enable : in  STD_LOGIC;
				  write_enable : in  STD_LOGIC;
				  ppn_in : in  STD_LOGIC_VECTOR (3 downto 0);
				  page_offset : in  STD_LOGIC_VECTOR (6 downto 0);
				  data_bus_in : in  PAGE;
				  clk : in  STD_LOGIC;
				  ppn_out : out STD_LOGIC_VECTOR (3 downto 0);
				  data_bus_out : out  STD_LOGIC_VECTOR (31 downto 0));
	end component;
	
	component PageTable is
		 Port ( read_enable : in  STD_LOGIC;
				  write_enable : in  STD_LOGIC;
				  vpn : in  STD_LOGIC_VECTOR (8 downto 0);
				  ppn_in : in  STD_LOGIC_VECTOR (3 downto 0); -- incoming ppn from MainMemory
				  clk : in  STD_LOGIC;
				  ppn_out : out  STD_LOGIC_VECTOR (3 downto 0); -- outgoing ppn to TLB
				  hit : out  STD_LOGIC);
	end component;
	
	component TLB is
		 Port ( read_enable : in  STD_LOGIC;
				  write_enable : in  STD_LOGIC;
				  vpn : in  STD_LOGIC_VECTOR (8 downto 0);
				  data_bus_in : in  STD_LOGIC_VECTOR (3 downto 0); -- input ppn
				  clk : in  STD_LOGIC;
				  data_bus_out : out  STD_LOGIC_VECTOR (3 downto 0); -- output ppn
				  hit : out  STD_LOGIC);
	end component;
	
	-- =========================================================================
	-- Signals:
	
	-- control signals
	SIGNAL tlb_read_en : STD_LOGIC := '0';
	SIGNAL tlb_write_en : STD_LOGIC := '0';
	SIGNAL tlb_hit : STD_LOGIC := '0';
	SIGNAL pt_read_en : STD_LOGIC := '0';
	SIGNAL pt_write_en : STD_LOGIC := '0';
	SIGNAL pt_hit : STD_LOGIC := '0';
	SIGNAL ram_read_en : STD_LOGIC := '0';
	SIGNAL ram_write_en : STD_LOGIC := '0';
	SIGNAL cache_read_en : STD_LOGIC := '0';
	SIGNAL cache_write_en : STD_LOGIC := '0';
	SIGNAL cache_hit : STD_LOGIC := '0';
	
	-- VA created generated by processor
	SIGNAL virtual_address : STD_LOGIC_VECTOR (15 downto 0); 
	ALIAS vpn : STD_LOGIC_VECTOR(8 downto 0) is virtual_address(15 downto 7);
	ALIAS page_offset : STD_LOGIC_VECTOR(6 downto 0) is virtual_address(6 downto 0);
	
	-- ppn signals
	SIGNAL ppn_out_tlb : STD_LOGIC_VECTOR(3 downto 0);
	SIGNAL ppn_out_pt : STD_LOGIC_VECTOR(3 downto 0);
	SIGNAL ppn_out_ram : STD_LOGIC_VECTOR(3 downto 0);
	
	-- data signals
	SIGNAL cache_data_out : STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL ram_data_out : STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL disk_data_out : PAGE;
	
	-- cache block address
	SIGNAL cache_block_address : STD_LOGIC_VECTOR(10 downto 0);
	
	-- =========================================================================
	-- Enumerated type declaration and state signal declaration
   SIGNAL State : state_type := Init;

	-- =========================================================================
	-- array of VAs and index
	TYPE data10in16 is ARRAY(0 to 9) of STD_LOGIC_VECTOR(15 downto 0);
	SIGNAL VA_memory : data10in16 := 
					("0100100110110101","1011101000111111","0000010011001011","0100110000001101",
					"0010101100010001","1101011010001111","1101100001011011","0011000100010000",
					"1011000010010010","0011011100101111");
	SIGNAL index : INTEGER RANGE 0 to 9;
	-- =========================================================================

begin

	DetermineState : Process(clk) is
	begin
		case State is
			when Init =>
				State <= Processor_State;
			--------------------
			when Processor_State =>
				State <= TLB_Read;
			--------------------
			when Cache_Read =>
				if (cache_hit = '1') then
					State <= Processor_State;
				else
					State <= RAM_Read;
				end if;
			--------------------
			when TLB_Read => 
				if (tlb_hit = '1') then
					State <= Cache_Read;
				else
					State <= PT_Read;
				end if;
			--------------------
			when PT_Read => 
				if (pt_hit = '1') then
					State <= TLB_Write;
				else
					State <= Disk_State;
				end if;
			--------------------
			when RAM_Read => 
				State <= Cache_Write;
			--------------------
			when Disk_State => 
				State <= RAM_Write;
			--------------------
			when Cache_Write => 
				State <= Cache_Read;
			--------------------
			when RAM_Write => 
				State <= PT_Write;
			--------------------
			when PT_Write => 
				State <= PT_Read;
			--------------------
			when TLB_Write => 
				State <= TLB_Read;
			--------------------
		end case;
	end Process;
	
	LogicProcess : Process(State) is
	begin
		case State is
			when Init =>
			-- setting all control signals.
				tlb_read_en <= '0';
				tlb_write_en <= '0';
				tlb_hit <= '0';
				pt_read_en <= '0';
				pt_write_en <= '0';
				pt_hit <= '0';
				ram_read_en <= '0';
				ram_write_en <= '0';
				cache_read_en <= '0';
				cache_write_en <= '0';
				cache_hit <= '0';
				
			when Processor_State =>
			-- setting all control signals.
				tlb_read_en <= '0';
				tlb_write_en <= '0';
				tlb_hit <= '0';
				pt_read_en <= '0';
				pt_write_en <= '0';
				pt_hit <= '0';
				ram_read_en <= '0';
				ram_write_en <= '0';
				cache_read_en <= '0';
				cache_write_en <= '0';
				cache_hit <= '0';
				
				virtual_address <= (others => '0');
				ppn_out_tlb <= (others => '0');
				ppn_out_pt <= (others => '0');
				ppn_out_ram <= (others => '0');
				cache_data_out <= (others => '0');
				ram_data_out <= (others => '0');
				disk_data_out <= (others => (others => '0'));
				cache_block_address <= (others => '0');
				
				virtual_address <= VA_memory(index);
				index <= index + 1;
			----------------------------------------
			when Cache_Read =>
				-- setting all control signals.
				tlb_read_en <= '0';
				tlb_write_en <= '0';
				tlb_hit <= '0';
				pt_read_en <= '0';
				pt_write_en <= '0';
				pt_hit <= '0';
				ram_read_en <= '0';
				ram_write_en <= '0';
				cache_read_en <= '1';
				cache_write_en <= '0';
				cache_hit <= '0';
				
			----------------------------------------
			when TLB_Read => 
				tlb_read_en <= '1';
				tlb_write_en <= '0';
				tlb_hit <= '0';
				pt_read_en <= '0';
				pt_write_en <= '0';
				pt_hit <= '0';
				ram_read_en <= '0';
				ram_write_en <= '0';
				cache_read_en <= '0';
				cache_write_en <= '0';
				cache_hit <= '0';
				
			----------------------------------------
			when PT_Read => 
				tlb_read_en <= '0';
				tlb_write_en <= '0';
				tlb_hit <= '0';
				pt_read_en <= '1';
				pt_write_en <= '0';
				pt_hit <= '0';
				ram_read_en <= '0';
				ram_write_en <= '0';
				cache_read_en <= '0';
				cache_write_en <= '0';
				cache_hit <= '0';
				
				cache_block_address <= ppn_out_tlb & page_offset;
			----------------------------------------
			when RAM_Read => 
				tlb_read_en <= '0';
				tlb_write_en <= '0';
				tlb_hit <= '0';
				pt_read_en <= '0';
				pt_write_en <= '0';
				pt_hit <= '0';
				ram_read_en <= '1';
				ram_write_en <= '0';
				cache_read_en <= '0';
				cache_write_en <= '0';
				cache_hit <= '0';
				
			----------------------------------------
			when Disk_State => 
				tlb_read_en <= '0';
				tlb_write_en <= '0';
				tlb_hit <= '0';
				pt_read_en <= '0';
				pt_write_en <= '0';
				pt_hit <= '0';
				ram_read_en <= '0';
				ram_write_en <= '0';
				cache_read_en <= '0';
				cache_write_en <= '0';
				cache_hit <= '0';
				
			----------------------------------------
			when Cache_Write => 
				tlb_read_en <= '0';
				tlb_write_en <= '0';
				tlb_hit <= '0';
				pt_read_en <= '0';
				pt_write_en <= '0';
				pt_hit <= '0';
				ram_read_en <= '0';
				ram_write_en <= '0';
				cache_read_en <= '0';
				cache_write_en <= '1';
				cache_hit <= '0';
				
			----------------------------------------
			when RAM_Write => 
				tlb_read_en <= '0';
				tlb_write_en <= '0';
				tlb_hit <= '0';
				pt_read_en <= '0';
				pt_write_en <= '0';
				pt_hit <= '0';
				ram_read_en <= '0';
				ram_write_en <= '1';
				cache_read_en <= '0';
				cache_write_en <= '0';
				cache_hit <= '0';
				
			----------------------------------------
			when PT_Write => 
				tlb_read_en <= '0';
				tlb_write_en <= '0';
				tlb_hit <= '0';
				pt_read_en <= '0';
				pt_write_en <= '1';
				pt_hit <= '0';
				ram_read_en <= '0';
				ram_write_en <= '0';
				cache_read_en <= '0';
				cache_write_en <= '0';
				cache_hit <= '0';
				
			----------------------------------------
			when TLB_Write => 
				tlb_read_en <= '0';
				tlb_write_en <= '1';
				tlb_hit <= '0';
				pt_read_en <= '0';
				pt_write_en <= '0';
				pt_hit <= '0';
				ram_read_en <= '0';
				ram_write_en <= '0';
				cache_read_en <= '0';
				cache_write_en <= '0';
				cache_hit <= '0';
				
			----------------------------------------
		end case;
	end Process;
	
	state_out_Process: Process(clk) is
	begin
		state_out <= State;
	end Process;
	
	data_out_Process : Process(State) is
	begin
		if (state = Cache_Read) then
			data_out <= cache_data_out;
		end if;
	end Process;
	
	Cache_Component : Cache(TwoWaySetAssociative) PORT MAP ( cache_read_en, cache_write_en, cache_block_address, 
												  ram_data_out, clk, cache_hit, cache_data_out );
	
	TLB_Component : TLB(FullAssociative) PORT MAP ( tlb_read_en, tlb_write_en, vpn, ppn_out_pt,
											 clk, ppn_out_tlb, tlb_hit);
	
	PT_Component : PageTable PORT MAP ( pt_read_en, pt_write_en, vpn, ppn_out_ram,
													clk, ppn_out_pt, pt_hit);
	
	RAM_Component : MainMemory PORT MAP ( ram_read_en, ram_write_en, ppn_out_pt, page_offset,
													  disk_data_out, clk, ppn_out_ram, ram_data_out);
													  
end Behavioral;

