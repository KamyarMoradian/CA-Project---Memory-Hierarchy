library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
library work;
    use work.Types.ALL;

entity Processor is
    Port ( clk : in  STD_LOGIC;
           tlb_v : in  STD_LOGIC;
           cache_v : in  STD_LOGIC;
			  state_out : out state_type;
           data_out : out  STD_LOGIC_VECTOR (31 downto 0));
end Processor;

architecture Behavioral of Processor is

	-- =========================================================================
	-- Signals:
	
	-- control signals
	SIGNAL tlb_v0_read_en : STD_LOGIC := '0';
	SIGNAL tlb_v0_write_en : STD_LOGIC := '0';
	SIGNAL tlb_v0_hit : STD_LOGIC := '0';
	SIGNAL tlb_v1_read_en : STD_LOGIC := '0';
	SIGNAL tlb_v1_write_en : STD_LOGIC := '0';
	SIGNAL tlb_v1_hit : STD_LOGIC := '0';
	SIGNAL tlb_hit : STD_LOGIC := '0';
	SIGNAL pt_read_en : STD_LOGIC := '0';
	SIGNAL pt_write_en : STD_LOGIC := '0';
	SIGNAL pt_hit : STD_LOGIC := '0';
	SIGNAL ram_read_en : STD_LOGIC := '0';
	SIGNAL ram_write_en : STD_LOGIC := '0';
	SIGNAL disc_read_en : STD_LOGIC := '0';
	SIGNAL cache_v0_read_en : STD_LOGIC := '0';
	SIGNAL cache_v0_write_en : STD_LOGIC := '0';
	SIGNAL cache_v0_hit : STD_LOGIC := '0';
	SIGNAL cache_v1_read_en : STD_LOGIC := '0';
	SIGNAL cache_v1_write_en : STD_LOGIC := '0';
	SIGNAL cache_v1_hit : STD_LOGIC := '0';
	SIGNAL cache_hit : STD_LOGIC := '0';
	
	-- VA created generated by processor
	SIGNAL virtual_address : STD_LOGIC_VECTOR (15 downto 0); 
	ALIAS vpn : STD_LOGIC_VECTOR(8 downto 0) is virtual_address(15 downto 7);
	ALIAS page_offset : STD_LOGIC_VECTOR(6 downto 0) is virtual_address(6 downto 0);
	
	-- ppn signals
	SIGNAL ppn_v0_out_tlb : STD_LOGIC_VECTOR(3 downto 0);
	SIGNAL ppn_v1_out_tlb : STD_LOGIC_VECTOR(3 downto 0);
	SIGNAL ppn_out_tlb : STD_LOGIC_VECTOR(3 downto 0);
	SIGNAL ppn_out_pt : STD_LOGIC_VECTOR(3 downto 0);
	SIGNAL ppn_out_ram : STD_LOGIC_VECTOR(3 downto 0);
	
	-- data signals
	SIGNAL cache_v0_data_out : STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL cache_v1_data_out : STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL ram_data_out : STD_LOGIC_VECTOR(63 downto 0);
	SIGNAL disc_data_out : PAGE;
	
	-- cache block address
	SIGNAL cache_v0_block_address : STD_LOGIC_VECTOR(10 downto 0);
	SIGNAL cache_v1_block_address : STD_LOGIC_VECTOR(10 downto 0);
	
	-- ram clock
	SIGNAL ram_clk : INTEGER;
	-- =========================================================================
	-- Enumerated type declaration and state signal declaration
   SIGNAL present_state : state_type := Init;
   SIGNAL next_state : state_type;

	-- =========================================================================
	-- array of VAs and index
	TYPE data14in16 is ARRAY(0 to 13) of STD_LOGIC_VECTOR(15 downto 0);
	SIGNAL VA_memory : data14in16 := 
					("0000000000000000","0000000000000100","0000000000001000","0000000000001100",
					"0000000000010000","0000000000000000","0000000000000100","0000000000001000",
					"0000000000001100","0000000000010000","0010000000000000","0010000000000100",
					"0010000000001000","0010000000001100");
--					,"1101100001011000","1101100001011100",
--					"1101100001100000","1101100001100100","0000000000000100","0000000000001000",
--					"0000000000001100","0000000000010000"
	SIGNAL index : INTEGER RANGE 0 to 14;
	
	-- =========================================================================

begin
	DeterminePresentState : Process(clk) is
	begin
		if (clk'event) then
			present_state <= next_state after 50 ns;
		end if;
	end Process;

	DetermineState : Process(clk) is
	begin
		if (present_state'STABLE AND FALLING_EDGE(clk)) then
			case present_state is
				when Init =>
					next_state <= Processor_State;
					
				--------------------
				when Processor_State =>
					next_state <= TLB_Read;
				--------------------
				when Cache_Read =>
					if (cache_hit = '1') then
						next_state <= Processor_State;
					else
						next_state <= RAM_Read;
					end if;
				--------------------
				when TLB_Read => 
					if (tlb_hit = '1') then
						next_state <= Cache_Read;
						if (cache_v = '0') then
							cache_v0_block_address <= ppn_out_tlb & page_offset;
						else
							cache_v1_block_address <= ppn_out_tlb & page_offset;
						end if;
					else
						next_state <= PT_Read;
					end if;
				--------------------
				when PT_Read => 
					if (pt_hit = '1') then
						next_state <= TLB_Write;
					else
						next_state <= Disc_State;
					end if;
				--------------------
				when RAM_Read => 
					next_state <= Cache_Write;
					
				--------------------
				when Disc_State =>
					next_state <= RAM_Write;
				--------------------
				when Cache_Write => 
					next_state <= Cache_Read;
				--------------------
				when RAM_Write =>
					next_state <= PT_Write;
				--------------------
				when PT_Write => 
					next_state <= PT_Read;
				--------------------
				when TLB_Write => 
					next_state <= TLB_Read;
				--------------------
			end case;
		end if;
	end Process;
	
	LogicProcess : Process(present_state) is
	begin
		tlb_v0_read_en <= '0';
		tlb_v1_read_en <= '0';
		tlb_v0_write_en <= '0';
		tlb_v1_write_en <= '0';
		pt_read_en <= '0';
		pt_write_en <= '0';
		ram_read_en <= '0';
		cache_v0_read_en <= '0';
		cache_v1_read_en <= '0';
		cache_v0_write_en <= '0';
		cache_v1_write_en <= '0';
		disc_read_en <= '0';
	
		case present_state is
			when Processor_State =>
				virtual_address <= VA_memory(index);
				if (cache_v = '0') then
					data_out <= cache_v0_data_out;
				else
					data_out <= cache_v1_data_out;
				end if;
				index <= (index + 1) mod 14;
			----------------------------------------
			when Cache_Read =>
				if (cache_v = '0') then
					cache_v0_read_en <= '1';
				else 
					cache_v1_read_en <= '1';
				end if;
			----------------------------------------
			when TLB_Read => 
				if (tlb_v = '0') then
					tlb_v0_read_en <= '1';
				else
					tlb_v1_read_en <= '1';
				end if;

			----------------------------------------
			when PT_Read => 
				pt_read_en <= '1';
				
			----------------------------------------
			when RAM_Read => 
				ram_read_en <= '1';

			----------------------------------------
			when Disc_State => 
				disc_read_en <= '1';

			----------------------------------------
			when Cache_Write => 
				if (cache_v = '0') then
					cache_v0_write_en <= '1';
				else
					cache_v1_write_en <= '1';
				end if;

			----------------------------------------
			when PT_Write => 
				pt_write_en <= '1';

			----------------------------------------
			when TLB_Write => 
				if (tlb_v = '0') then
					tlb_v0_write_en <= '1';
				else
					tlb_v1_write_en <= '1';
				end if;

			----------------------------------------
			when others =>
				null;
		end case;
	end Process;
	
	state_out_Process: Process(present_state) is
	begin
		state_out <= present_state;
	end Process;
	
	ram_clk_Process : Process(clk) is
	begin
		if (present_state = RAM_Write AND ram_clk >= 2) then
			ram_write_en <= '1';
		else 
			ram_write_en <= '0';
		end if;
		if (present_state = RAM_Write) then
			ram_clk <= (ram_clk + 1) mod 5;
		else ram_clk <= 0;
		end if;
	end Process;
	
	cache_hit_process : Process (cache_v0_hit, cache_v1_hit) is
	begin
		if (cache_v = '0') then
			cache_hit <= cache_v0_hit;
		else
			cache_hit <= cache_v1_hit;
		end if;
	end Process;
	
	tlb_hit_process : Process (tlb_v0_hit, tlb_v1_hit) is
	begin
		if (tlb_v = '0') then
			tlb_hit <= tlb_v0_hit;
		else
			tlb_hit <= tlb_v1_hit;
		end if;
	end Process;
	
	ppn_out_tlb_process : Process (ppn_v0_out_tlb, ppn_v1_out_tlb) is
	begin
		if (tlb_v = '0') then
			ppn_out_tlb <= ppn_v0_out_tlb;
		else
			ppn_out_tlb <= ppn_v1_out_tlb;
		end if;
	end Process;
	
	Cache_v0_Component : entity work.Cache(DirectMapped) PORT MAP 
												 ( cache_v0_read_en, cache_v0_write_en, cache_v0_block_address, 
												   ram_data_out, clk, cache_v0_hit, cache_v0_data_out );
	Cache_v1_Component : entity work.Cache(TwoWaySetAssociative) PORT MAP 
												 ( cache_v1_read_en, cache_v1_write_en, cache_v1_block_address, 
												   ram_data_out, clk, cache_v1_hit, cache_v1_data_out );
	
	TLB_v0_Component : entity work.TLB(FullAssociative) PORT MAP 
											( tlb_v0_read_en, tlb_v0_write_en, vpn, ppn_out_pt,
											  clk, ppn_v0_out_tlb, tlb_v0_hit);
	TLB_v1_Component : entity work.TLB(FourWaySetAssociative) PORT MAP 
											( tlb_v1_read_en, tlb_v1_write_en, vpn, ppn_out_pt,
											  clk, ppn_v1_out_tlb, tlb_v1_hit);
	
	PT_Component : entity work.PageTable PORT MAP ( pt_read_en, pt_write_en, vpn, ppn_out_ram,
																	clk, ppn_out_pt, pt_hit);
	
	RAM_Component : entity work.MainMemory PORT MAP ( ram_read_en, ram_write_en, ppn_out_pt, page_offset,
																	  disc_data_out, clk, ppn_out_ram, ram_data_out);
	
	Disc_Component : entity work.HardDisc PORT MAP ( disc_read_en, clk, vpn, disc_data_out);
	
end Behavioral;

